// <Student_ID> <Name>

// e.g. 110123456 王大明
// Add your ID and name to FIRST line of file, or you will get 5 points penalty
module exam1_B(
    input wire clk,
    input wire rst,
    output reg [15:0] out// You can modify "reg" to "wire" if needed
);
    //Your design here

endmodule

// You can add any module you need.
// Make sure you include all modules you used in this problem.